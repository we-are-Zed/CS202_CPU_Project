    module setchar(
        input clk,
        input rst,
        
    );
    
    endmodule