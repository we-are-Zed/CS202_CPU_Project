module  seg_transform 
(
input [15:0]seg_in,
output [31:0]seg_out
);
wire [3:0]seg_in1,seg_in2,seg_in3,seg_in4;
assign seg_in1=seg_in[3:0];
assign seg_in2=seg_in[7:4];
assign seg_in3=seg_in[11:8];
assign seg_in4=seg_in[15:12];
//输入的数据，分为4段，每一段对应一个数码管输出
reg [7:0]seg1,seg2,seg3,seg4;
assign seg_out={seg4,seg3,seg2,seg1};
always@* begin
case(seg_in1)
4'b0000: seg1 <= 8'b11000000;  //  0
            4'b0001: seg1 <= 8'b11111001;  //  1
            4'b0010: seg1 <= 8'b10100100;  //  2
            4'b0011: seg1 <= 8'b10110000;  //  3
            4'b0100: seg1 <= 8'b10011001;  //  4
            4'b0101: seg1 <= 8'b10010010;  //  5
            4'b0110: seg1 <= 8'b10000010;  //  6
            4'b0111: seg1 <= 8'b11111000;  //  7
            4'b1000: seg1 <= 8'b10000000;  //  8
            4'b1001: seg1 <= 8'b10010000;  //  9
            4'b1010: seg1 <= 8'b10001000;  //  A
            4'b1011: seg1 <= 8'b10000011;  //  b
            4'b1100: seg1 <= 8'b11000110;  //  C
            4'b1101: seg1 <= 8'b10100001;  //  d
            4'b1110: seg1 <= 8'b10000110;  //  E
            4'b1111: seg1 <= 8'b11111111;  //  F  
            default: seg1 <= 8'b00000000;
endcase
end
always@* begin
case(seg_in2)
4'b0000: seg2 <= 8'b11000000;  //  0
            4'b0001: seg2 <= 8'b11111001;  //  1
            4'b0010: seg2 <= 8'b10100100;  //  2
            4'b0011: seg2 <= 8'b10110000;  //  3
            4'b0100: seg2 <= 8'b10011001;  //  4
            4'b0101: seg2 <= 8'b10010010;  //  5
            4'b0110: seg2 <= 8'b10000010;  //  6
            4'b0111: seg2 <= 8'b11111000;  //  7
            4'b1000: seg2 <= 8'b10000000;  //  8
            4'b1001: seg2 <= 8'b10010000;  //  9
            4'b1010: seg2 <= 8'b10001000;  //  A
            4'b1011: seg2 <= 8'b10000011;  //  b
            4'b1100: seg2 <= 8'b11000110;  //  C
            4'b1101: seg2 <= 8'b10100001;  //  d
            4'b1110: seg2 <= 8'b10000110;  //  E
            4'b1111: seg2 <= 8'b11111111;  //  F  
            default: seg2 <= 8'b00000000;
endcase
end
always@ *begin
case(seg_in3)
4'b0000: seg3 <= 8'b11000000;  //  0
            4'b0001: seg3 <= 8'b11111001;  //  1
            4'b0010: seg3 <= 8'b10100100;  //  2
            4'b0011: seg3 <= 8'b10110000;  //  3
            4'b0100: seg3 <= 8'b10011001;  //  4
            4'b0101: seg3 <= 8'b10010010;  //  5
            4'b0110: seg3 <= 8'b10000010;  //  6
            4'b0111: seg3 <= 8'b11111000;  //  7
            4'b1000: seg3 <= 8'b10000000;  //  8
            4'b1001: seg3 <= 8'b10010000;  //  9
            4'b1010: seg3 <= 8'b10001000;  //  A
            4'b1011: seg3 <= 8'b10000011;  //  b
            4'b1100: seg3 <= 8'b11000110;  //  C
            4'b1101: seg3 <= 8'b10100001;  //  d
            4'b1110: seg3 <= 8'b10000110;  //  E
            4'b1111: seg3 <= 8'b11111111;  //  F  
            default: seg3 <= 8'b00000000;
endcase
end
always@ *begin
case(seg_in4)
4'b0000: seg4 <= 8'b11000000;  //  0
            4'b0001: seg4 <= 8'b11111001;  //  1
            4'b0010: seg4 <= 8'b10100100;  //  2
            4'b0011: seg4 <= 8'b10110000;  //  3
            4'b0100: seg4 <= 8'b10011001;  //  4
            4'b0101: seg4 <= 8'b10010010;  //  5
            4'b0110: seg4 <= 8'b10000010;  //  6
            4'b0111: seg4 <= 8'b11111000;  //  7
            4'b1000: seg4 <= 8'b10000000;  //  8
            4'b1001: seg4 <= 8'b10010000;  //  9
            4'b1010: seg4 <= 8'b10001000;  //  A
            4'b1011: seg4 <= 8'b10000011;  //  b
            4'b1100: seg4 <= 8'b11000110;  //  C
            4'b1101: seg4 <= 8'b10100001;  //  d
            4'b1110: seg4 <= 8'b10000110;  //  E
            4'b1111: seg4 <= 8'b11111111;  //  F  
            default: seg1 <= 8'b00000000;
endcase
end


endmodule